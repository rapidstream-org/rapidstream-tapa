endmodule  // {{ module.name }}
